library IEEE;
use IEEE.std_logic_1164.all;


entity gc_cntr is
  port (
    reset : in  std_logic;    -- Async. active-high reset.
    clk   : in  std_logic;    -- Rising-edge-active clock.
	 ena : std_logic;
    q     : out std_logic_vector(7 downto 0) -- Counter output.
    );
end entity;


architecture arch of gc_cntr is
  signal cntr_r, cntr_x : std_logic_vector(7 downto 0); -- Current and next counter state.
begin

  -- Compute next counter state from current counter state.
  with cntr_r select cntr_x(0) <= not cntr_r(0) when "00000000",
                                  not cntr_r(0) when "00000011",
                                  not cntr_r(0) when "00000110",
                                  not cntr_r(0) when "00000101",
                                  not cntr_r(0) when "00001100",
                                  not cntr_r(0) when "00001111",
                                  not cntr_r(0) when "00001010",
                                  not cntr_r(0) when "00001001",
                                  not cntr_r(0) when "00011000",
                                  not cntr_r(0) when "00011011",
                                  not cntr_r(0) when "00011110",
                                  not cntr_r(0) when "00011101",
                                  not cntr_r(0) when "00010100",
                                  not cntr_r(0) when "00010111",
                                  not cntr_r(0) when "00010010",
                                  not cntr_r(0) when "00010001",
                                  not cntr_r(0) when "00110000",
                                  not cntr_r(0) when "00110011",
                                  not cntr_r(0) when "00110110",
                                  not cntr_r(0) when "00110101",
                                  not cntr_r(0) when "00111100",
                                  not cntr_r(0) when "00111111",
                                  not cntr_r(0) when "00111010",
                                  not cntr_r(0) when "00111001",
                                  not cntr_r(0) when "00101000",
                                  not cntr_r(0) when "00101011",
                                  not cntr_r(0) when "00101110",
                                  not cntr_r(0) when "00101101",
                                  not cntr_r(0) when "00100100",
                                  not cntr_r(0) when "00100111",
                                  not cntr_r(0) when "00100010",
                                  not cntr_r(0) when "00100001",
                                  not cntr_r(0) when "01100000",
                                  not cntr_r(0) when "01100011",
                                  not cntr_r(0) when "01100110",
                                  not cntr_r(0) when "01100101",
                                  not cntr_r(0) when "01101100",
                                  not cntr_r(0) when "01101111",
                                  not cntr_r(0) when "01101010",
                                  not cntr_r(0) when "01101001",
                                  not cntr_r(0) when "01111000",
                                  not cntr_r(0) when "01111011",
                                  not cntr_r(0) when "01111110",
                                  not cntr_r(0) when "01111101",
                                  not cntr_r(0) when "01110100",
                                  not cntr_r(0) when "01110111",
                                  not cntr_r(0) when "01110010",
                                  not cntr_r(0) when "01110001",
                                  not cntr_r(0) when "01010000",
                                  not cntr_r(0) when "01010011",
                                  not cntr_r(0) when "01010110",
                                  not cntr_r(0) when "01010101",
                                  not cntr_r(0) when "01011100",
                                  not cntr_r(0) when "01011111",
                                  not cntr_r(0) when "01011010",
                                  not cntr_r(0) when "01011001",
                                  not cntr_r(0) when "01001000",
                                  not cntr_r(0) when "01001011",
                                  not cntr_r(0) when "01001110",
                                  not cntr_r(0) when "01001101",
                                  not cntr_r(0) when "01000100",
                                  not cntr_r(0) when "01000111",
                                  not cntr_r(0) when "01000010",
                                  not cntr_r(0) when "01000001",
                                  not cntr_r(0) when "11000000",
                                  not cntr_r(0) when "11000011",
                                  not cntr_r(0) when "11000110",
                                  not cntr_r(0) when "11000101",
                                  not cntr_r(0) when "11001100",
                                  not cntr_r(0) when "11001111",
                                  not cntr_r(0) when "11001010",
                                  not cntr_r(0) when "11001001",
                                  not cntr_r(0) when "11011000",
                                  not cntr_r(0) when "11011011",
                                  not cntr_r(0) when "11011110",
                                  not cntr_r(0) when "11011101",
                                  not cntr_r(0) when "11010100",
                                  not cntr_r(0) when "11010111",
                                  not cntr_r(0) when "11010010",
                                  not cntr_r(0) when "11010001",
                                  not cntr_r(0) when "11110000",
                                  not cntr_r(0) when "11110011",
                                  not cntr_r(0) when "11110110",
                                  not cntr_r(0) when "11110101",
                                  not cntr_r(0) when "11111100",
                                  not cntr_r(0) when "11111111",
                                  not cntr_r(0) when "11111010",
                                  not cntr_r(0) when "11111001",
                                  not cntr_r(0) when "11101000",
                                  not cntr_r(0) when "11101011",
                                  not cntr_r(0) when "11101110",
                                  not cntr_r(0) when "11101101",
                                  not cntr_r(0) when "11100100",
                                  not cntr_r(0) when "11100111",
                                  not cntr_r(0) when "11100010",
                                  not cntr_r(0) when "11100001",
                                  not cntr_r(0) when "10100000",
                                  not cntr_r(0) when "10100011",
                                  not cntr_r(0) when "10100110",
                                  not cntr_r(0) when "10100101",
                                  not cntr_r(0) when "10101100",
                                  not cntr_r(0) when "10101111",
                                  not cntr_r(0) when "10101010",
                                  not cntr_r(0) when "10101001",
                                  not cntr_r(0) when "10111000",
                                  not cntr_r(0) when "10111011",
                                  not cntr_r(0) when "10111110",
                                  not cntr_r(0) when "10111101",
                                  not cntr_r(0) when "10110100",
                                  not cntr_r(0) when "10110111",
                                  not cntr_r(0) when "10110010",
                                  not cntr_r(0) when "10110001",
                                  not cntr_r(0) when "10010000",
                                  not cntr_r(0) when "10010011",
                                  not cntr_r(0) when "10010110",
                                  not cntr_r(0) when "10010101",
                                  not cntr_r(0) when "10011100",
                                  not cntr_r(0) when "10011111",
                                  not cntr_r(0) when "10011010",
                                  not cntr_r(0) when "10011001",
                                  not cntr_r(0) when "10001000",
                                  not cntr_r(0) when "10001011",
                                  not cntr_r(0) when "10001110",
                                  not cntr_r(0) when "10001101",
                                  not cntr_r(0) when "10000100",
                                  not cntr_r(0) when "10000111",
                                  not cntr_r(0) when "10000010",
                                  not cntr_r(0) when "10000001",
                                      cntr_r(0) when others;
  with cntr_r select cntr_x(1) <= not cntr_r(1) when "00000001",
                                  not cntr_r(1) when "00000111",
                                  not cntr_r(1) when "00001101",
                                  not cntr_r(1) when "00001011",
                                  not cntr_r(1) when "00011001",
                                  not cntr_r(1) when "00011111",
                                  not cntr_r(1) when "00010101",
                                  not cntr_r(1) when "00010011",
                                  not cntr_r(1) when "00110001",
                                  not cntr_r(1) when "00110111",
                                  not cntr_r(1) when "00111101",
                                  not cntr_r(1) when "00111011",
                                  not cntr_r(1) when "00101001",
                                  not cntr_r(1) when "00101111",
                                  not cntr_r(1) when "00100101",
                                  not cntr_r(1) when "00100011",
                                  not cntr_r(1) when "01100001",
                                  not cntr_r(1) when "01100111",
                                  not cntr_r(1) when "01101101",
                                  not cntr_r(1) when "01101011",
                                  not cntr_r(1) when "01111001",
                                  not cntr_r(1) when "01111111",
                                  not cntr_r(1) when "01110101",
                                  not cntr_r(1) when "01110011",
                                  not cntr_r(1) when "01010001",
                                  not cntr_r(1) when "01010111",
                                  not cntr_r(1) when "01011101",
                                  not cntr_r(1) when "01011011",
                                  not cntr_r(1) when "01001001",
                                  not cntr_r(1) when "01001111",
                                  not cntr_r(1) when "01000101",
                                  not cntr_r(1) when "01000011",
                                  not cntr_r(1) when "11000001",
                                  not cntr_r(1) when "11000111",
                                  not cntr_r(1) when "11001101",
                                  not cntr_r(1) when "11001011",
                                  not cntr_r(1) when "11011001",
                                  not cntr_r(1) when "11011111",
                                  not cntr_r(1) when "11010101",
                                  not cntr_r(1) when "11010011",
                                  not cntr_r(1) when "11110001",
                                  not cntr_r(1) when "11110111",
                                  not cntr_r(1) when "11111101",
                                  not cntr_r(1) when "11111011",
                                  not cntr_r(1) when "11101001",
                                  not cntr_r(1) when "11101111",
                                  not cntr_r(1) when "11100101",
                                  not cntr_r(1) when "11100011",
                                  not cntr_r(1) when "10100001",
                                  not cntr_r(1) when "10100111",
                                  not cntr_r(1) when "10101101",
                                  not cntr_r(1) when "10101011",
                                  not cntr_r(1) when "10111001",
                                  not cntr_r(1) when "10111111",
                                  not cntr_r(1) when "10110101",
                                  not cntr_r(1) when "10110011",
                                  not cntr_r(1) when "10010001",
                                  not cntr_r(1) when "10010111",
                                  not cntr_r(1) when "10011101",
                                  not cntr_r(1) when "10011011",
                                  not cntr_r(1) when "10001001",
                                  not cntr_r(1) when "10001111",
                                  not cntr_r(1) when "10000101",
                                  not cntr_r(1) when "10000011",
                                      cntr_r(1) when others;
  with cntr_r select cntr_x(2) <= not cntr_r(2) when "00000010",
                                  not cntr_r(2) when "00001110",
                                  not cntr_r(2) when "00011010",
                                  not cntr_r(2) when "00010110",
                                  not cntr_r(2) when "00110010",
                                  not cntr_r(2) when "00111110",
                                  not cntr_r(2) when "00101010",
                                  not cntr_r(2) when "00100110",
                                  not cntr_r(2) when "01100010",
                                  not cntr_r(2) when "01101110",
                                  not cntr_r(2) when "01111010",
                                  not cntr_r(2) when "01110110",
                                  not cntr_r(2) when "01010010",
                                  not cntr_r(2) when "01011110",
                                  not cntr_r(2) when "01001010",
                                  not cntr_r(2) when "01000110",
                                  not cntr_r(2) when "11000010",
                                  not cntr_r(2) when "11001110",
                                  not cntr_r(2) when "11011010",
                                  not cntr_r(2) when "11010110",
                                  not cntr_r(2) when "11110010",
                                  not cntr_r(2) when "11111110",
                                  not cntr_r(2) when "11101010",
                                  not cntr_r(2) when "11100110",
                                  not cntr_r(2) when "10100010",
                                  not cntr_r(2) when "10101110",
                                  not cntr_r(2) when "10111010",
                                  not cntr_r(2) when "10110110",
                                  not cntr_r(2) when "10010010",
                                  not cntr_r(2) when "10011110",
                                  not cntr_r(2) when "10001010",
                                  not cntr_r(2) when "10000110",
                                      cntr_r(2) when others;
  with cntr_r select cntr_x(3) <= not cntr_r(3) when "00000100",
                                  not cntr_r(3) when "00011100",
                                  not cntr_r(3) when "00110100",
                                  not cntr_r(3) when "00101100",
                                  not cntr_r(3) when "01100100",
                                  not cntr_r(3) when "01111100",
                                  not cntr_r(3) when "01010100",
                                  not cntr_r(3) when "01001100",
                                  not cntr_r(3) when "11000100",
                                  not cntr_r(3) when "11011100",
                                  not cntr_r(3) when "11110100",
                                  not cntr_r(3) when "11101100",
                                  not cntr_r(3) when "10100100",
                                  not cntr_r(3) when "10111100",
                                  not cntr_r(3) when "10010100",
                                  not cntr_r(3) when "10001100",
                                      cntr_r(3) when others;
  with cntr_r select cntr_x(4) <= not cntr_r(4) when "00001000",
                                  not cntr_r(4) when "00111000",
                                  not cntr_r(4) when "01101000",
                                  not cntr_r(4) when "01011000",
                                  not cntr_r(4) when "11001000",
                                  not cntr_r(4) when "11111000",
                                  not cntr_r(4) when "10101000",
                                  not cntr_r(4) when "10011000",
                                      cntr_r(4) when others;
  with cntr_r select cntr_x(5) <= not cntr_r(5) when "00010000",
                                  not cntr_r(5) when "01110000",
                                  not cntr_r(5) when "11010000",
                                  not cntr_r(5) when "10110000",
                                      cntr_r(5) when others;
  with cntr_r select cntr_x(6) <= not cntr_r(6) when "00100000",
                                  not cntr_r(6) when "11100000",
                                      cntr_r(6) when others;
  with cntr_r select cntr_x(7) <= not cntr_r(7) when "01000000",
                                  not cntr_r(7) when "10000000",
                                      cntr_r(7) when others;

  process(reset,clk)
  begin
    if reset = '1' then
      cntr_r <= "00000000"; -- Reset counter value.
    elsif rising_edge(clk) then
		if ena = '1' then
			cntr_r <= cntr_x; -- Update counter value.
		end if;
    end if;
  end process;

  q <= cntr_r; -- Output counter value.

end architecture;
